
// file: ibert_ultrascale_gth_0.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_ibert_ultrascale_gth_0
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module example_ibert_ultrascale_gth_0
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////

`define C_NUM_GTH_QUADS 4
`define C_GTH_REFCLKS_USED 4
module example_ibert_ultrascale_gth_0
(
  // GT top level ports
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txn_o,
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txp_o,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]    	gth_rxn_i,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]   	gth_rxp_i,
  input                           	gth_sysclkp_i,
  input                           	gth_sysclkn_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0n_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1n_i,
  output kus_dl_sel,
  output fpga_sel_18,
  output rst_clks_18_b,
  input ccb_hardrst_b,
  input ccb_soft_rst,
  input done,
  output RX12_I2C_ENA, 
  output RX12_CS_B,
  output RX12_RST_B,
  output TX12_I2C_ENA,
  output TX12_CS_B,
  output TX12_RST_B,
  output B04_I2C_ENA,
  output B04_CS_B,
  output B04_RST_B,
  output DAQ_SPY_SEL_18,
  input B04_INT_B,
  input B04_PRESENT_B
);

  //
  // Ibert refclk internal signals
  //
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk1_i;        	
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk11_i; 
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk1_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_1_i;
  wire                        gth_sysclk_i;


  //
  // Refclk IBUFDS instantiations
  //
    IBUFDS_GTE3 u_buf_gth_q0_clk0
      (
        .O            (gth_refclk0_i[0]),
        .ODIV2        (gth_odiv2_0_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[0]),
        .IB           (gth_refclk0n_i[0])
      );

    IBUFDS_GTE3 u_buf_gth_q0_clk1
      (
        .O            (gth_refclk1_i[0]),
        .ODIV2        (gth_odiv2_1_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[0]),
        .IB           (gth_refclk1n_i[0])
      );
    IBUFDS_GTE3 u_buf_gth_q1_clk0
      (
        .O            (gth_refclk0_i[1]),
        .ODIV2        (gth_odiv2_0_i[1]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[1]),
        .IB           (gth_refclk0n_i[1])
      );

    IBUFDS_GTE3 u_buf_gth_q1_clk1
      (
        .O            (gth_refclk1_i[1]),
        .ODIV2        (gth_odiv2_1_i[1]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[1]),
        .IB           (gth_refclk1n_i[1])
      );
    IBUFDS_GTE3 u_buf_gth_q2_clk0
      (
        .O            (gth_refclk0_i[2]),
        .ODIV2        (gth_odiv2_0_i[2]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[2]),
        .IB           (gth_refclk0n_i[2])
      );

    IBUFDS_GTE3 u_buf_gth_q2_clk1
      (
        .O            (gth_refclk1_i[2]),
        .ODIV2        (gth_odiv2_1_i[2]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[2]),
        .IB           (gth_refclk1n_i[2])
      );
    IBUFDS_GTE3 u_buf_gth_q3_clk0
      (
        .O            (gth_refclk0_i[3]),
        .ODIV2        (gth_odiv2_0_i[3]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[3]),
        .IB           (gth_refclk0n_i[3])
      );

    IBUFDS_GTE3 u_buf_gth_q3_clk1
      (
        .O            (gth_refclk1_i[3]),
        .ODIV2        (gth_odiv2_1_i[3]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[3]),
        .IB           (gth_refclk1n_i[3])
      );

  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gth_qrefclk0_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk1_i[0] = gth_refclk1_i[0];
  assign gth_qnorthrefclk0_i[0] = 1'b0;
  assign gth_qnorthrefclk1_i[0] = 1'b0;
  assign gth_qsouthrefclk0_i[0] = 1'b0;
  assign gth_qsouthrefclk1_i[0] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[0] = 1'b0;
  assign gth_qrefclk10_i[0] = 1'b0;
  assign gth_qrefclk01_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk11_i[0] = gth_refclk1_i[0];  
  assign gth_qnorthrefclk00_i[0] = 1'b0;
  assign gth_qnorthrefclk10_i[0] = 1'b0;
  assign gth_qnorthrefclk01_i[0] = 1'b0;
  assign gth_qnorthrefclk11_i[0] = 1'b0;  
  assign gth_qsouthrefclk00_i[0] = 1'b0;
  assign gth_qsouthrefclk10_i[0] = 1'b0;  
  assign gth_qsouthrefclk01_i[0] = 1'b0;
  assign gth_qsouthrefclk11_i[0] = 1'b0;

  assign gth_qrefclk0_i[1] = gth_refclk0_i[1];
  assign gth_qrefclk1_i[1] = gth_refclk1_i[1];
  assign gth_qnorthrefclk0_i[1] = 1'b0;
  assign gth_qnorthrefclk1_i[1] = 1'b0;
  assign gth_qsouthrefclk0_i[1] = 1'b0;
  assign gth_qsouthrefclk1_i[1] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[1] = 1'b0;
  assign gth_qrefclk10_i[1] = 1'b0;
  assign gth_qrefclk01_i[1] = gth_refclk0_i[1];
  assign gth_qrefclk11_i[1] = gth_refclk1_i[1];  
  assign gth_qnorthrefclk00_i[1] = 1'b0;
  assign gth_qnorthrefclk10_i[1] = 1'b0;
  assign gth_qnorthrefclk01_i[1] = 1'b0;
  assign gth_qnorthrefclk11_i[1] = 1'b0;  
  assign gth_qsouthrefclk00_i[1] = 1'b0;
  assign gth_qsouthrefclk10_i[1] = 1'b0;  
  assign gth_qsouthrefclk01_i[1] = 1'b0;
  assign gth_qsouthrefclk11_i[1] = 1'b0;

  assign gth_qrefclk0_i[2] = gth_refclk0_i[2];
  assign gth_qrefclk1_i[2] = gth_refclk1_i[2];
  assign gth_qnorthrefclk0_i[2] = 1'b0;
  assign gth_qnorthrefclk1_i[2] = 1'b0;
  assign gth_qsouthrefclk0_i[2] = 1'b0;
  assign gth_qsouthrefclk1_i[2] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[2] = 1'b0;
  assign gth_qrefclk10_i[2] = 1'b0;
  assign gth_qrefclk01_i[2] = gth_refclk0_i[2];
  assign gth_qrefclk11_i[2] = gth_refclk1_i[2];  
  assign gth_qnorthrefclk00_i[2] = 1'b0;
  assign gth_qnorthrefclk10_i[2] = 1'b0;
  assign gth_qnorthrefclk01_i[2] = 1'b0;
  assign gth_qnorthrefclk11_i[2] = 1'b0;  
  assign gth_qsouthrefclk00_i[2] = 1'b0;
  assign gth_qsouthrefclk10_i[2] = 1'b0;  
  assign gth_qsouthrefclk01_i[2] = 1'b0;
  assign gth_qsouthrefclk11_i[2] = 1'b0;

  assign gth_qrefclk0_i[3] = gth_refclk0_i[3];
  assign gth_qrefclk1_i[3] = gth_refclk1_i[3];
  assign gth_qnorthrefclk0_i[3] = 1'b0;
  assign gth_qnorthrefclk1_i[3] = 1'b0;
  assign gth_qsouthrefclk0_i[3] = 1'b0;
  assign gth_qsouthrefclk1_i[3] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[3] = 1'b0;
  assign gth_qrefclk10_i[3] = 1'b0;
  assign gth_qrefclk01_i[3] = gth_refclk0_i[3];
  assign gth_qrefclk11_i[3] = gth_refclk1_i[3];  
  assign gth_qnorthrefclk00_i[3] = 1'b0;
  assign gth_qnorthrefclk10_i[3] = 1'b0;
  assign gth_qnorthrefclk01_i[3] = 1'b0;
  assign gth_qnorthrefclk11_i[3] = 1'b0;  
  assign gth_qsouthrefclk00_i[3] = 1'b0;
  assign gth_qsouthrefclk10_i[3] = 1'b0;  
  assign gth_qsouthrefclk01_i[3] = 1'b0;
  assign gth_qsouthrefclk11_i[3] = 1'b0;

  assign kus_dl_sel    = 1'b1;
  assign fpga_sel_18   = 1'b0;
  assign rst_clks_18_b = 1'b1;
  assign RX12_I2C_ENA  = 1'b0;
  assign RX12_CS_B     = 1'b1;
  assign RX12_RST_B    = 1'b1;
  assign TX12_I2C_ENA  = 1'b0;
  assign TX12_CS_B     = 1'b1;
  assign TX12_RST_B    = 1'b1;
  assign B04_I2C_ENA   = 1'b0;
  assign B04_CS_B      = 1'b1;
  assign B04_RST_B     = 1'b1;

  //
  // Sysclock IBUFDS instantiation
  //
  IBUFGDS 
   #(.DIFF_TERM("FALSE"))
   u_ibufgds
    (
      .I(gth_sysclkp_i),
      .IB(gth_sysclkn_i),
      .O(gth_sysclk_i)
    );


  //
  // IBERT core instantiation
  //
  ibert_ultrascale_gth_0 u_ibert_gth_core
    (
      .txn_o(gth_txn_o),
      .txp_o(gth_txp_o),
      .rxn_i(gth_rxn_i),
      .rxp_i(gth_rxp_i),
      .clk(gth_sysclk_i),
      .gtrefclk0_i(gth_qrefclk0_i),
      .gtrefclk1_i(gth_qrefclk1_i),
      .gtnorthrefclk0_i(gth_qnorthrefclk0_i),
      .gtnorthrefclk1_i(gth_qnorthrefclk1_i),
      .gtsouthrefclk0_i(gth_qsouthrefclk0_i),
      .gtsouthrefclk1_i(gth_qsouthrefclk1_i),
      .gtrefclk00_i(gth_qrefclk00_i),
      .gtrefclk10_i(gth_qrefclk10_i),
      .gtrefclk01_i(gth_qrefclk01_i),
      .gtrefclk11_i(gth_qrefclk11_i),
      .gtnorthrefclk00_i(gth_qnorthrefclk00_i),
      .gtnorthrefclk10_i(gth_qnorthrefclk10_i),
      .gtnorthrefclk01_i(gth_qnorthrefclk01_i),
      .gtnorthrefclk11_i(gth_qnorthrefclk11_i),
      .gtsouthrefclk00_i(gth_qsouthrefclk00_i),
      .gtsouthrefclk10_i(gth_qsouthrefclk10_i),
      .gtsouthrefclk01_i(gth_qsouthrefclk01_i),
      .gtsouthrefclk11_i(gth_qsouthrefclk11_i)
    );

  vio_0 spy
    (
       .clk(gth_sysclk_i),
       .probe_out0(DAQ_SPY_SEL_18)
    );


endmodule
